`define version_major_cvi_ciris    4'd0
`define version_minor_cvi_ciris    6'd0
`define version_revision_cvi_ciris 22'd0